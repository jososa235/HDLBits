//problem found at: https://hdlbits.01xz.net/wiki/Sim/circuit1


module top_module (
    input a,
    input b,
    output q );//

    assign q = a & b; // Fix me

endmodule